module ALU()

reg[3:0] ALUControl;
always @(*)
    case(ALUOp)
    

    endcase

endmodule